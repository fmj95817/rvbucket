`ifndef BOOT_ROM_SVH
`define BOOT_ROM_SVH

`define BOOT_ROM_WORD_AW 5

`endif
