../../../sim/rtl/model/rom.sv