../../../sim/rtl/model/sram.sv