`ifndef BOOT_ROM_SVH
`define BOOT_ROM_SVH

`define BOOT_ROM_AW 4

`endif
