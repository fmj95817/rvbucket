module lsu(
    input           clk,
    input           rst_n,
    ldst_if.slave   ldst_src,
    ldst_if.master  ldst_gen
);
    assign ldst_gen.req_vld = ldst_src.req_vld;
    assign ldst_gen.req_pkt = ldst_src.req_pkt;
    assign ldst_src.req_rdy = ldst_gen.req_rdy;

    assign ldst_src.rsp_vld = ldst_gen.rsp_vld;
    assign ldst_src.rsp_pkt = ldst_gen.rsp_pkt;
    assign ldst_gen.rsp_rdy = ldst_src.rsp_rdy;
endmodule